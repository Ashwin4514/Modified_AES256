module decryptRound(in,key,out,thresholdVal);
input [127:0] in;
output [127:0] out;
input [127:0] key;
input [127:0] thresholdVal;
wire [127:0] SBO;
wire [127:0] SBRO;

inverseShiftRows r(in,SBRO);
inverseSubBytes s(SBRO,SBO,thresholdVal);
addRoundKey b(SBO,out,key);

endmodule