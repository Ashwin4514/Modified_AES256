module decryptor_tb;

reg [127:0] in;
wire [127:0] out;
reg [255:0] key;
reg [255:0] sbox_seed;

decryption c(in,key,out,sbox_seed);


initial begin

in=128'hc21bd6808b2e6508def33538894c31b2;
key=256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f;
sbox_seed=256'h000102030405060708090a0b0c0d0e0f101112131415161718191a1b1c1d1e1f;
$monitor("Inside Decryptor Testbench: in256= %h, key256= %h ,out256= %h",in,key,out);
//temp= 'h3205442b026d1e7773450f4f513877464e7f6a40191235257f6a2a6b64237c563b046c532c6c5f1f786f541062491f6e5227126b2a164b240b00597c754b246f632c056454146249200b65212363370e68247e004027754c25046a3d0b764c330d4d2d18653e0a5f1e09143710785f38796940116a4f1d5d3634054e331e7736357c1f167b542270601f0a5f382370603a7a4439126b391e5e4534643d1c0c4c260d473e256555187161327d494b18714b226c4511014e1d0d5a4568654c1d76553571314d0d664b197243250a3722070c5759187f68246469597c6335257e41;

end

endmodule